// Code your design here
`include "sfp.v"
// Code your testbench here
// or browse Examples
`include "sfp_tb.v"